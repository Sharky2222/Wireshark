-- Wire_Shark.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Wire_Shark is
	port (
		clk_clk                                   : in  std_logic                    := '0';             --                             clk.clk
		eth_tse_0_mac_mdio_connection_mdc         : out std_logic;                                       --   eth_tse_0_mac_mdio_connection.mdc
		eth_tse_0_mac_mdio_connection_mdio_in     : in  std_logic                    := '0';             --                                .mdio_in
		eth_tse_0_mac_mdio_connection_mdio_out    : out std_logic;                                       --                                .mdio_out
		eth_tse_0_mac_mdio_connection_mdio_oen    : out std_logic;                                       --                                .mdio_oen
		eth_tse_0_mac_rgmii_connection_rgmii_in   : in  std_logic_vector(3 downto 0) := (others => '0'); --  eth_tse_0_mac_rgmii_connection.rgmii_in
		eth_tse_0_mac_rgmii_connection_rgmii_out  : out std_logic_vector(3 downto 0);                    --                                .rgmii_out
		eth_tse_0_mac_rgmii_connection_rx_control : in  std_logic                    := '0';             --                                .rx_control
		eth_tse_0_mac_rgmii_connection_tx_control : out std_logic;                                       --                                .tx_control
		eth_tse_0_mac_status_connection_set_10    : in  std_logic                    := '0';             -- eth_tse_0_mac_status_connection.set_10
		eth_tse_0_mac_status_connection_set_1000  : in  std_logic                    := '0';             --                                .set_1000
		eth_tse_0_mac_status_connection_eth_mode  : out std_logic;                                       --                                .eth_mode
		eth_tse_0_mac_status_connection_ena_10    : out std_logic                                        --                                .ena_10
	);
end entity Wire_Shark;

architecture rtl of Wire_Shark is
	component PacketFilter is
		port (
			outData       : out std_logic_vector(31 downto 0);                    -- readdata
			inData        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			address       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			readTo        : in  std_logic                     := 'X';             -- read
			writeTo       : in  std_logic                     := 'X';             -- write
			avsChannel    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			startofpacket : in  std_logic                     := 'X';             -- startofpacket
			endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clock         : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X'              -- reset
		);
	end component PacketFilter;

	component Wire_Shark_SGDMA_RX is
		port (
			clk                           : in  std_logic                     := 'X';             -- clk
			system_reset_n                : in  std_logic                     := 'X';             -- reset_n
			csr_chipselect                : in  std_logic                     := 'X';             -- chipselect
			csr_address                   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			csr_read                      : in  std_logic                     := 'X';             -- read
			csr_write                     : in  std_logic                     := 'X';             -- write
			csr_writedata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			csr_readdata                  : out std_logic_vector(31 downto 0);                    -- readdata
			descriptor_read_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			descriptor_read_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			descriptor_read_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			descriptor_read_address       : out std_logic_vector(31 downto 0);                    -- address
			descriptor_read_read          : out std_logic;                                        -- read
			descriptor_write_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			descriptor_write_address      : out std_logic_vector(31 downto 0);                    -- address
			descriptor_write_write        : out std_logic;                                        -- write
			descriptor_write_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			csr_irq                       : out std_logic;                                        -- irq
			in_startofpacket              : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket                : in  std_logic                     := 'X';             -- endofpacket
			in_data                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_valid                      : in  std_logic                     := 'X';             -- valid
			in_ready                      : out std_logic;                                        -- ready
			in_empty                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			in_error                      : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- error
			m_write_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			m_write_address               : out std_logic_vector(31 downto 0);                    -- address
			m_write_write                 : out std_logic;                                        -- write
			m_write_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			m_write_byteenable            : out std_logic_vector(3 downto 0)                      -- byteenable
		);
	end component Wire_Shark_SGDMA_RX;

	component Wire_Shark_SGDMA_TX is
		port (
			clk                           : in  std_logic                     := 'X';             -- clk
			system_reset_n                : in  std_logic                     := 'X';             -- reset_n
			csr_chipselect                : in  std_logic                     := 'X';             -- chipselect
			csr_address                   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			csr_read                      : in  std_logic                     := 'X';             -- read
			csr_write                     : in  std_logic                     := 'X';             -- write
			csr_writedata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			csr_readdata                  : out std_logic_vector(31 downto 0);                    -- readdata
			descriptor_read_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			descriptor_read_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			descriptor_read_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			descriptor_read_address       : out std_logic_vector(31 downto 0);                    -- address
			descriptor_read_read          : out std_logic;                                        -- read
			descriptor_write_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			descriptor_write_address      : out std_logic_vector(31 downto 0);                    -- address
			descriptor_write_write        : out std_logic;                                        -- write
			descriptor_write_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			csr_irq                       : out std_logic;                                        -- irq
			m_read_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m_read_readdatavalid          : in  std_logic                     := 'X';             -- readdatavalid
			m_read_waitrequest            : in  std_logic                     := 'X';             -- waitrequest
			m_read_address                : out std_logic_vector(31 downto 0);                    -- address
			m_read_read                   : out std_logic;                                        -- read
			out_data                      : out std_logic_vector(31 downto 0);                    -- data
			out_valid                     : out std_logic;                                        -- valid
			out_ready                     : in  std_logic                     := 'X';             -- ready
			out_endofpacket               : out std_logic;                                        -- endofpacket
			out_startofpacket             : out std_logic;                                        -- startofpacket
			out_empty                     : out std_logic_vector(1 downto 0);                     -- empty
			out_error                     : out std_logic                                         -- error
		);
	end component Wire_Shark_SGDMA_TX;

	component Wire_Shark_TSE_MAC is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			reg_addr      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			reg_data_out  : out std_logic_vector(31 downto 0);                    -- readdata
			reg_rd        : in  std_logic                     := 'X';             -- read
			reg_data_in   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			reg_wr        : in  std_logic                     := 'X';             -- write
			reg_busy      : out std_logic;                                        -- waitrequest
			tx_clk        : in  std_logic                     := 'X';             -- clk
			rx_clk        : in  std_logic                     := 'X';             -- clk
			set_10        : in  std_logic                     := 'X';             -- set_10
			set_1000      : in  std_logic                     := 'X';             -- set_1000
			eth_mode      : out std_logic;                                        -- eth_mode
			ena_10        : out std_logic;                                        -- ena_10
			rgmii_in      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- rgmii_in
			rgmii_out     : out std_logic_vector(3 downto 0);                     -- rgmii_out
			rx_control    : in  std_logic                     := 'X';             -- rx_control
			tx_control    : out std_logic;                                        -- tx_control
			ff_rx_clk     : in  std_logic                     := 'X';             -- clk
			ff_tx_clk     : in  std_logic                     := 'X';             -- clk
			ff_rx_data    : out std_logic_vector(31 downto 0);                    -- data
			ff_rx_eop     : out std_logic;                                        -- endofpacket
			rx_err        : out std_logic_vector(5 downto 0);                     -- error
			ff_rx_mod     : out std_logic_vector(1 downto 0);                     -- empty
			ff_rx_rdy     : in  std_logic                     := 'X';             -- ready
			ff_rx_sop     : out std_logic;                                        -- startofpacket
			ff_rx_dval    : out std_logic;                                        -- valid
			ff_tx_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			ff_tx_eop     : in  std_logic                     := 'X';             -- endofpacket
			ff_tx_err     : in  std_logic                     := 'X';             -- error
			ff_tx_mod     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			ff_tx_rdy     : out std_logic;                                        -- ready
			ff_tx_sop     : in  std_logic                     := 'X';             -- startofpacket
			ff_tx_wren    : in  std_logic                     := 'X';             -- valid
			mdc           : out std_logic;                                        -- mdc
			mdio_in       : in  std_logic                     := 'X';             -- mdio_in
			mdio_out      : out std_logic;                                        -- mdio_out
			mdio_oen      : out std_logic;                                        -- mdio_oen
			magic_wakeup  : out std_logic;                                        -- magic_wakeup
			magic_sleep_n : in  std_logic                     := 'X';             -- magic_sleep_n
			ff_tx_crc_fwd : in  std_logic                     := 'X';             -- ff_tx_crc_fwd
			ff_tx_septy   : out std_logic;                                        -- ff_tx_septy
			tx_ff_uflow   : out std_logic;                                        -- tx_ff_uflow
			ff_tx_a_full  : out std_logic;                                        -- ff_tx_a_full
			ff_tx_a_empty : out std_logic;                                        -- ff_tx_a_empty
			rx_err_stat   : out std_logic_vector(17 downto 0);                    -- rx_err_stat
			rx_frm_type   : out std_logic_vector(3 downto 0);                     -- rx_frm_type
			ff_rx_dsav    : out std_logic;                                        -- ff_rx_dsav
			ff_rx_a_full  : out std_logic;                                        -- ff_rx_a_full
			ff_rx_a_empty : out std_logic                                         -- ff_rx_a_empty
		);
	end component Wire_Shark_TSE_MAC;

	component Wire_Shark_UART is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component Wire_Shark_UART;

	component Wire_Shark_demultiplexer_0 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset_n            : in  std_logic                     := 'X';             -- reset_n
			in_data            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_valid           : in  std_logic                     := 'X';             -- valid
			in_ready           : out std_logic;                                        -- ready
			in_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			in_empty           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			in_channel         : in  std_logic                     := 'X';             -- channel
			out0_data          : out std_logic_vector(31 downto 0);                    -- data
			out0_valid         : out std_logic;                                        -- valid
			out0_ready         : in  std_logic                     := 'X';             -- ready
			out0_startofpacket : out std_logic;                                        -- startofpacket
			out0_endofpacket   : out std_logic;                                        -- endofpacket
			out0_empty         : out std_logic_vector(1 downto 0);                     -- empty
			out1_data          : out std_logic_vector(31 downto 0);                    -- data
			out1_valid         : out std_logic;                                        -- valid
			out1_ready         : in  std_logic                     := 'X';             -- ready
			out1_startofpacket : out std_logic;                                        -- startofpacket
			out1_endofpacket   : out std_logic;                                        -- endofpacket
			out1_empty         : out std_logic_vector(1 downto 0)                      -- empty
		);
	end component Wire_Shark_demultiplexer_0;

	component Wire_Shark_descriptor_memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component Wire_Shark_descriptor_memory;

	component Wire_Shark_nios2e is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(15 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(15 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component Wire_Shark_nios2e;

	component Wire_Shark_onchip_memory_nios is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component Wire_Shark_onchip_memory_nios;

	component Wire_Shark_pll_0 is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component Wire_Shark_pll_0;

	component Wire_Shark_mm_interconnect_0 is
		port (
			clk_0_clk_clk                            : in  std_logic                     := 'X';             -- clk
			nios2e_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2e_data_master_address               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			nios2e_data_master_waitrequest           : out std_logic;                                        -- waitrequest
			nios2e_data_master_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2e_data_master_read                  : in  std_logic                     := 'X';             -- read
			nios2e_data_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			nios2e_data_master_write                 : in  std_logic                     := 'X';             -- write
			nios2e_data_master_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2e_data_master_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			nios2e_instruction_master_address        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			nios2e_instruction_master_waitrequest    : out std_logic;                                        -- waitrequest
			nios2e_instruction_master_read           : in  std_logic                     := 'X';             -- read
			nios2e_instruction_master_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			SGDMA_RX_descriptor_read_address         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			SGDMA_RX_descriptor_read_waitrequest     : out std_logic;                                        -- waitrequest
			SGDMA_RX_descriptor_read_read            : in  std_logic                     := 'X';             -- read
			SGDMA_RX_descriptor_read_readdata        : out std_logic_vector(31 downto 0);                    -- readdata
			SGDMA_RX_descriptor_read_readdatavalid   : out std_logic;                                        -- readdatavalid
			SGDMA_RX_descriptor_write_address        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			SGDMA_RX_descriptor_write_waitrequest    : out std_logic;                                        -- waitrequest
			SGDMA_RX_descriptor_write_write          : in  std_logic                     := 'X';             -- write
			SGDMA_RX_descriptor_write_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			SGDMA_RX_m_write_address                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			SGDMA_RX_m_write_waitrequest             : out std_logic;                                        -- waitrequest
			SGDMA_RX_m_write_byteenable              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			SGDMA_RX_m_write_write                   : in  std_logic                     := 'X';             -- write
			SGDMA_RX_m_write_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			SGDMA_TX_descriptor_read_address         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			SGDMA_TX_descriptor_read_waitrequest     : out std_logic;                                        -- waitrequest
			SGDMA_TX_descriptor_read_read            : in  std_logic                     := 'X';             -- read
			SGDMA_TX_descriptor_read_readdata        : out std_logic_vector(31 downto 0);                    -- readdata
			SGDMA_TX_descriptor_read_readdatavalid   : out std_logic;                                        -- readdatavalid
			SGDMA_TX_descriptor_write_address        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			SGDMA_TX_descriptor_write_waitrequest    : out std_logic;                                        -- waitrequest
			SGDMA_TX_descriptor_write_write          : in  std_logic                     := 'X';             -- write
			SGDMA_TX_descriptor_write_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			SGDMA_TX_m_read_address                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			SGDMA_TX_m_read_waitrequest              : out std_logic;                                        -- waitrequest
			SGDMA_TX_m_read_read                     : in  std_logic                     := 'X';             -- read
			SGDMA_TX_m_read_readdata                 : out std_logic_vector(31 downto 0);                    -- readdata
			SGDMA_TX_m_read_readdatavalid            : out std_logic;                                        -- readdatavalid
			descriptor_memory_s1_address             : out std_logic_vector(9 downto 0);                     -- address
			descriptor_memory_s1_write               : out std_logic;                                        -- write
			descriptor_memory_s1_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			descriptor_memory_s1_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			descriptor_memory_s1_byteenable          : out std_logic_vector(3 downto 0);                     -- byteenable
			descriptor_memory_s1_chipselect          : out std_logic;                                        -- chipselect
			descriptor_memory_s1_clken               : out std_logic;                                        -- clken
			Filter_0_avalon_slave_0_address          : out std_logic_vector(3 downto 0);                     -- address
			Filter_0_avalon_slave_0_write            : out std_logic;                                        -- write
			Filter_0_avalon_slave_0_read             : out std_logic;                                        -- read
			Filter_0_avalon_slave_0_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Filter_0_avalon_slave_0_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			Filter_0_avalon_slave_0_chipselect       : out std_logic;                                        -- chipselect
			nios2e_debug_mem_slave_address           : out std_logic_vector(8 downto 0);                     -- address
			nios2e_debug_mem_slave_write             : out std_logic;                                        -- write
			nios2e_debug_mem_slave_read              : out std_logic;                                        -- read
			nios2e_debug_mem_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2e_debug_mem_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			nios2e_debug_mem_slave_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2e_debug_mem_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			nios2e_debug_mem_slave_debugaccess       : out std_logic;                                        -- debugaccess
			onchip_memory_nios_s1_address            : out std_logic_vector(11 downto 0);                    -- address
			onchip_memory_nios_s1_write              : out std_logic;                                        -- write
			onchip_memory_nios_s1_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory_nios_s1_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory_nios_s1_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory_nios_s1_chipselect         : out std_logic;                                        -- chipselect
			onchip_memory_nios_s1_clken              : out std_logic;                                        -- clken
			SGDMA_RX_csr_address                     : out std_logic_vector(3 downto 0);                     -- address
			SGDMA_RX_csr_write                       : out std_logic;                                        -- write
			SGDMA_RX_csr_read                        : out std_logic;                                        -- read
			SGDMA_RX_csr_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			SGDMA_RX_csr_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			SGDMA_RX_csr_chipselect                  : out std_logic;                                        -- chipselect
			SGDMA_TX_csr_address                     : out std_logic_vector(3 downto 0);                     -- address
			SGDMA_TX_csr_write                       : out std_logic;                                        -- write
			SGDMA_TX_csr_read                        : out std_logic;                                        -- read
			SGDMA_TX_csr_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			SGDMA_TX_csr_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			SGDMA_TX_csr_chipselect                  : out std_logic;                                        -- chipselect
			TSE_MAC_control_port_address             : out std_logic_vector(7 downto 0);                     -- address
			TSE_MAC_control_port_write               : out std_logic;                                        -- write
			TSE_MAC_control_port_read                : out std_logic;                                        -- read
			TSE_MAC_control_port_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			TSE_MAC_control_port_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			TSE_MAC_control_port_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			UART_avalon_jtag_slave_address           : out std_logic_vector(0 downto 0);                     -- address
			UART_avalon_jtag_slave_write             : out std_logic;                                        -- write
			UART_avalon_jtag_slave_read              : out std_logic;                                        -- read
			UART_avalon_jtag_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			UART_avalon_jtag_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			UART_avalon_jtag_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			UART_avalon_jtag_slave_chipselect        : out std_logic                                         -- chipselect
		);
	end component Wire_Shark_mm_interconnect_0;

	component Wire_Shark_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component Wire_Shark_irq_mapper;

	component Wire_Shark_avalon_st_adapter is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk        : in  std_logic                     := 'X';             -- clk
			in_rst_0_reset      : in  std_logic                     := 'X';             -- reset
			in_0_data           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_0_valid          : in  std_logic                     := 'X';             -- valid
			in_0_ready          : out std_logic;                                        -- ready
			in_0_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_0_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			in_0_empty          : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			out_0_data          : out std_logic_vector(31 downto 0);                    -- data
			out_0_valid         : out std_logic;                                        -- valid
			out_0_ready         : in  std_logic                     := 'X';             -- ready
			out_0_startofpacket : out std_logic;                                        -- startofpacket
			out_0_endofpacket   : out std_logic;                                        -- endofpacket
			out_0_empty         : out std_logic_vector(1 downto 0);                     -- empty
			out_0_error         : out std_logic_vector(5 downto 0)                      -- error
		);
	end component Wire_Shark_avalon_st_adapter;

	component Wire_Shark_avalon_st_adapter_001 is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk        : in  std_logic                     := 'X';             -- clk
			in_rst_0_reset      : in  std_logic                     := 'X';             -- reset
			in_0_data           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_0_valid          : in  std_logic                     := 'X';             -- valid
			in_0_ready          : out std_logic;                                        -- ready
			in_0_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_0_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			in_0_empty          : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			out_0_data          : out std_logic_vector(31 downto 0);                    -- data
			out_0_startofpacket : out std_logic;                                        -- startofpacket
			out_0_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component Wire_Shark_avalon_st_adapter_001;

	component Wire_Shark_avalon_st_adapter_002 is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk        : in  std_logic                     := 'X';             -- clk
			in_rst_0_reset      : in  std_logic                     := 'X';             -- reset
			in_0_data           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_0_valid          : in  std_logic                     := 'X';             -- valid
			in_0_ready          : out std_logic;                                        -- ready
			in_0_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_0_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			in_0_empty          : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			in_0_error          : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- error
			out_0_data          : out std_logic_vector(31 downto 0);                    -- data
			out_0_valid         : out std_logic;                                        -- valid
			out_0_ready         : in  std_logic                     := 'X';             -- ready
			out_0_startofpacket : out std_logic;                                        -- startofpacket
			out_0_endofpacket   : out std_logic;                                        -- endofpacket
			out_0_empty         : out std_logic_vector(1 downto 0);                     -- empty
			out_0_channel       : out std_logic                                         -- channel
		);
	end component Wire_Shark_avalon_st_adapter_002;

	component wire_shark_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component wire_shark_rst_controller;

	component wire_shark_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component wire_shark_rst_controller_001;

	signal sgdma_tx_out_valid                                       : std_logic;                     -- SGDMA_TX:out_valid -> TSE_MAC:ff_tx_wren
	signal sgdma_tx_out_data                                        : std_logic_vector(31 downto 0); -- SGDMA_TX:out_data -> TSE_MAC:ff_tx_data
	signal sgdma_tx_out_ready                                       : std_logic;                     -- TSE_MAC:ff_tx_rdy -> SGDMA_TX:out_ready
	signal sgdma_tx_out_startofpacket                               : std_logic;                     -- SGDMA_TX:out_startofpacket -> TSE_MAC:ff_tx_sop
	signal sgdma_tx_out_endofpacket                                 : std_logic;                     -- SGDMA_TX:out_endofpacket -> TSE_MAC:ff_tx_eop
	signal sgdma_tx_out_error                                       : std_logic;                     -- SGDMA_TX:out_error -> TSE_MAC:ff_tx_err
	signal sgdma_tx_out_empty                                       : std_logic_vector(1 downto 0);  -- SGDMA_TX:out_empty -> TSE_MAC:ff_tx_mod
	signal pll_0_outclk0_clk                                        : std_logic;                     -- pll_0:outclk_0 -> [TSE_MAC:rx_clk, TSE_MAC:tx_clk]
	signal nios2e_debug_reset_request_reset                         : std_logic;                     -- nios2e:debug_reset_request -> [pll_0:rst, rst_controller:reset_in0, rst_controller:reset_in1, rst_controller_001:reset_in0]
	signal nios2e_data_master_readdata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2e_data_master_readdata -> nios2e:d_readdata
	signal nios2e_data_master_waitrequest                           : std_logic;                     -- mm_interconnect_0:nios2e_data_master_waitrequest -> nios2e:d_waitrequest
	signal nios2e_data_master_debugaccess                           : std_logic;                     -- nios2e:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2e_data_master_debugaccess
	signal nios2e_data_master_address                               : std_logic_vector(15 downto 0); -- nios2e:d_address -> mm_interconnect_0:nios2e_data_master_address
	signal nios2e_data_master_byteenable                            : std_logic_vector(3 downto 0);  -- nios2e:d_byteenable -> mm_interconnect_0:nios2e_data_master_byteenable
	signal nios2e_data_master_read                                  : std_logic;                     -- nios2e:d_read -> mm_interconnect_0:nios2e_data_master_read
	signal nios2e_data_master_write                                 : std_logic;                     -- nios2e:d_write -> mm_interconnect_0:nios2e_data_master_write
	signal nios2e_data_master_writedata                             : std_logic_vector(31 downto 0); -- nios2e:d_writedata -> mm_interconnect_0:nios2e_data_master_writedata
	signal sgdma_tx_descriptor_read_readdata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:SGDMA_TX_descriptor_read_readdata -> SGDMA_TX:descriptor_read_readdata
	signal sgdma_tx_descriptor_read_waitrequest                     : std_logic;                     -- mm_interconnect_0:SGDMA_TX_descriptor_read_waitrequest -> SGDMA_TX:descriptor_read_waitrequest
	signal sgdma_tx_descriptor_read_address                         : std_logic_vector(31 downto 0); -- SGDMA_TX:descriptor_read_address -> mm_interconnect_0:SGDMA_TX_descriptor_read_address
	signal sgdma_tx_descriptor_read_read                            : std_logic;                     -- SGDMA_TX:descriptor_read_read -> mm_interconnect_0:SGDMA_TX_descriptor_read_read
	signal sgdma_tx_descriptor_read_readdatavalid                   : std_logic;                     -- mm_interconnect_0:SGDMA_TX_descriptor_read_readdatavalid -> SGDMA_TX:descriptor_read_readdatavalid
	signal sgdma_rx_descriptor_read_readdata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:SGDMA_RX_descriptor_read_readdata -> SGDMA_RX:descriptor_read_readdata
	signal sgdma_rx_descriptor_read_waitrequest                     : std_logic;                     -- mm_interconnect_0:SGDMA_RX_descriptor_read_waitrequest -> SGDMA_RX:descriptor_read_waitrequest
	signal sgdma_rx_descriptor_read_address                         : std_logic_vector(31 downto 0); -- SGDMA_RX:descriptor_read_address -> mm_interconnect_0:SGDMA_RX_descriptor_read_address
	signal sgdma_rx_descriptor_read_read                            : std_logic;                     -- SGDMA_RX:descriptor_read_read -> mm_interconnect_0:SGDMA_RX_descriptor_read_read
	signal sgdma_rx_descriptor_read_readdatavalid                   : std_logic;                     -- mm_interconnect_0:SGDMA_RX_descriptor_read_readdatavalid -> SGDMA_RX:descriptor_read_readdatavalid
	signal sgdma_tx_descriptor_write_waitrequest                    : std_logic;                     -- mm_interconnect_0:SGDMA_TX_descriptor_write_waitrequest -> SGDMA_TX:descriptor_write_waitrequest
	signal sgdma_tx_descriptor_write_address                        : std_logic_vector(31 downto 0); -- SGDMA_TX:descriptor_write_address -> mm_interconnect_0:SGDMA_TX_descriptor_write_address
	signal sgdma_tx_descriptor_write_write                          : std_logic;                     -- SGDMA_TX:descriptor_write_write -> mm_interconnect_0:SGDMA_TX_descriptor_write_write
	signal sgdma_tx_descriptor_write_writedata                      : std_logic_vector(31 downto 0); -- SGDMA_TX:descriptor_write_writedata -> mm_interconnect_0:SGDMA_TX_descriptor_write_writedata
	signal sgdma_rx_descriptor_write_waitrequest                    : std_logic;                     -- mm_interconnect_0:SGDMA_RX_descriptor_write_waitrequest -> SGDMA_RX:descriptor_write_waitrequest
	signal sgdma_rx_descriptor_write_address                        : std_logic_vector(31 downto 0); -- SGDMA_RX:descriptor_write_address -> mm_interconnect_0:SGDMA_RX_descriptor_write_address
	signal sgdma_rx_descriptor_write_write                          : std_logic;                     -- SGDMA_RX:descriptor_write_write -> mm_interconnect_0:SGDMA_RX_descriptor_write_write
	signal sgdma_rx_descriptor_write_writedata                      : std_logic_vector(31 downto 0); -- SGDMA_RX:descriptor_write_writedata -> mm_interconnect_0:SGDMA_RX_descriptor_write_writedata
	signal nios2e_instruction_master_readdata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2e_instruction_master_readdata -> nios2e:i_readdata
	signal nios2e_instruction_master_waitrequest                    : std_logic;                     -- mm_interconnect_0:nios2e_instruction_master_waitrequest -> nios2e:i_waitrequest
	signal nios2e_instruction_master_address                        : std_logic_vector(15 downto 0); -- nios2e:i_address -> mm_interconnect_0:nios2e_instruction_master_address
	signal nios2e_instruction_master_read                           : std_logic;                     -- nios2e:i_read -> mm_interconnect_0:nios2e_instruction_master_read
	signal sgdma_tx_m_read_readdata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:SGDMA_TX_m_read_readdata -> SGDMA_TX:m_read_readdata
	signal sgdma_tx_m_read_waitrequest                              : std_logic;                     -- mm_interconnect_0:SGDMA_TX_m_read_waitrequest -> SGDMA_TX:m_read_waitrequest
	signal sgdma_tx_m_read_address                                  : std_logic_vector(31 downto 0); -- SGDMA_TX:m_read_address -> mm_interconnect_0:SGDMA_TX_m_read_address
	signal sgdma_tx_m_read_read                                     : std_logic;                     -- SGDMA_TX:m_read_read -> mm_interconnect_0:SGDMA_TX_m_read_read
	signal sgdma_tx_m_read_readdatavalid                            : std_logic;                     -- mm_interconnect_0:SGDMA_TX_m_read_readdatavalid -> SGDMA_TX:m_read_readdatavalid
	signal sgdma_rx_m_write_waitrequest                             : std_logic;                     -- mm_interconnect_0:SGDMA_RX_m_write_waitrequest -> SGDMA_RX:m_write_waitrequest
	signal sgdma_rx_m_write_address                                 : std_logic_vector(31 downto 0); -- SGDMA_RX:m_write_address -> mm_interconnect_0:SGDMA_RX_m_write_address
	signal sgdma_rx_m_write_byteenable                              : std_logic_vector(3 downto 0);  -- SGDMA_RX:m_write_byteenable -> mm_interconnect_0:SGDMA_RX_m_write_byteenable
	signal sgdma_rx_m_write_write                                   : std_logic;                     -- SGDMA_RX:m_write_write -> mm_interconnect_0:SGDMA_RX_m_write_write
	signal sgdma_rx_m_write_writedata                               : std_logic_vector(31 downto 0); -- SGDMA_RX:m_write_writedata -> mm_interconnect_0:SGDMA_RX_m_write_writedata
	signal mm_interconnect_0_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:UART_avalon_jtag_slave_chipselect -> UART:av_chipselect
	signal mm_interconnect_0_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- UART:av_readdata -> mm_interconnect_0:UART_avalon_jtag_slave_readdata
	signal mm_interconnect_0_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- UART:av_waitrequest -> mm_interconnect_0:UART_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:UART_avalon_jtag_slave_address -> UART:av_address
	signal mm_interconnect_0_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:UART_avalon_jtag_slave_read -> mm_interconnect_0_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:UART_avalon_jtag_slave_write -> mm_interconnect_0_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:UART_avalon_jtag_slave_writedata -> UART:av_writedata
	signal mm_interconnect_0_filter_0_avalon_slave_0_chipselect     : std_logic;                     -- mm_interconnect_0:Filter_0_avalon_slave_0_chipselect -> Filter_0:chipselect
	signal mm_interconnect_0_filter_0_avalon_slave_0_readdata       : std_logic_vector(31 downto 0); -- Filter_0:outData -> mm_interconnect_0:Filter_0_avalon_slave_0_readdata
	signal mm_interconnect_0_filter_0_avalon_slave_0_address        : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Filter_0_avalon_slave_0_address -> Filter_0:address
	signal mm_interconnect_0_filter_0_avalon_slave_0_read           : std_logic;                     -- mm_interconnect_0:Filter_0_avalon_slave_0_read -> Filter_0:readTo
	signal mm_interconnect_0_filter_0_avalon_slave_0_write          : std_logic;                     -- mm_interconnect_0:Filter_0_avalon_slave_0_write -> Filter_0:writeTo
	signal mm_interconnect_0_filter_0_avalon_slave_0_writedata      : std_logic_vector(31 downto 0); -- mm_interconnect_0:Filter_0_avalon_slave_0_writedata -> Filter_0:inData
	signal mm_interconnect_0_tse_mac_control_port_readdata          : std_logic_vector(31 downto 0); -- TSE_MAC:reg_data_out -> mm_interconnect_0:TSE_MAC_control_port_readdata
	signal mm_interconnect_0_tse_mac_control_port_waitrequest       : std_logic;                     -- TSE_MAC:reg_busy -> mm_interconnect_0:TSE_MAC_control_port_waitrequest
	signal mm_interconnect_0_tse_mac_control_port_address           : std_logic_vector(7 downto 0);  -- mm_interconnect_0:TSE_MAC_control_port_address -> TSE_MAC:reg_addr
	signal mm_interconnect_0_tse_mac_control_port_read              : std_logic;                     -- mm_interconnect_0:TSE_MAC_control_port_read -> TSE_MAC:reg_rd
	signal mm_interconnect_0_tse_mac_control_port_write             : std_logic;                     -- mm_interconnect_0:TSE_MAC_control_port_write -> TSE_MAC:reg_wr
	signal mm_interconnect_0_tse_mac_control_port_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:TSE_MAC_control_port_writedata -> TSE_MAC:reg_data_in
	signal mm_interconnect_0_sgdma_rx_csr_chipselect                : std_logic;                     -- mm_interconnect_0:SGDMA_RX_csr_chipselect -> SGDMA_RX:csr_chipselect
	signal mm_interconnect_0_sgdma_rx_csr_readdata                  : std_logic_vector(31 downto 0); -- SGDMA_RX:csr_readdata -> mm_interconnect_0:SGDMA_RX_csr_readdata
	signal mm_interconnect_0_sgdma_rx_csr_address                   : std_logic_vector(3 downto 0);  -- mm_interconnect_0:SGDMA_RX_csr_address -> SGDMA_RX:csr_address
	signal mm_interconnect_0_sgdma_rx_csr_read                      : std_logic;                     -- mm_interconnect_0:SGDMA_RX_csr_read -> SGDMA_RX:csr_read
	signal mm_interconnect_0_sgdma_rx_csr_write                     : std_logic;                     -- mm_interconnect_0:SGDMA_RX_csr_write -> SGDMA_RX:csr_write
	signal mm_interconnect_0_sgdma_rx_csr_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:SGDMA_RX_csr_writedata -> SGDMA_RX:csr_writedata
	signal mm_interconnect_0_sgdma_tx_csr_chipselect                : std_logic;                     -- mm_interconnect_0:SGDMA_TX_csr_chipselect -> SGDMA_TX:csr_chipselect
	signal mm_interconnect_0_sgdma_tx_csr_readdata                  : std_logic_vector(31 downto 0); -- SGDMA_TX:csr_readdata -> mm_interconnect_0:SGDMA_TX_csr_readdata
	signal mm_interconnect_0_sgdma_tx_csr_address                   : std_logic_vector(3 downto 0);  -- mm_interconnect_0:SGDMA_TX_csr_address -> SGDMA_TX:csr_address
	signal mm_interconnect_0_sgdma_tx_csr_read                      : std_logic;                     -- mm_interconnect_0:SGDMA_TX_csr_read -> SGDMA_TX:csr_read
	signal mm_interconnect_0_sgdma_tx_csr_write                     : std_logic;                     -- mm_interconnect_0:SGDMA_TX_csr_write -> SGDMA_TX:csr_write
	signal mm_interconnect_0_sgdma_tx_csr_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:SGDMA_TX_csr_writedata -> SGDMA_TX:csr_writedata
	signal mm_interconnect_0_nios2e_debug_mem_slave_readdata        : std_logic_vector(31 downto 0); -- nios2e:debug_mem_slave_readdata -> mm_interconnect_0:nios2e_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2e_debug_mem_slave_waitrequest     : std_logic;                     -- nios2e:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2e_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2e_debug_mem_slave_debugaccess     : std_logic;                     -- mm_interconnect_0:nios2e_debug_mem_slave_debugaccess -> nios2e:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2e_debug_mem_slave_address         : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2e_debug_mem_slave_address -> nios2e:debug_mem_slave_address
	signal mm_interconnect_0_nios2e_debug_mem_slave_read            : std_logic;                     -- mm_interconnect_0:nios2e_debug_mem_slave_read -> nios2e:debug_mem_slave_read
	signal mm_interconnect_0_nios2e_debug_mem_slave_byteenable      : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2e_debug_mem_slave_byteenable -> nios2e:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2e_debug_mem_slave_write           : std_logic;                     -- mm_interconnect_0:nios2e_debug_mem_slave_write -> nios2e:debug_mem_slave_write
	signal mm_interconnect_0_nios2e_debug_mem_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2e_debug_mem_slave_writedata -> nios2e:debug_mem_slave_writedata
	signal mm_interconnect_0_onchip_memory_nios_s1_chipselect       : std_logic;                     -- mm_interconnect_0:onchip_memory_nios_s1_chipselect -> onchip_memory_nios:chipselect
	signal mm_interconnect_0_onchip_memory_nios_s1_readdata         : std_logic_vector(31 downto 0); -- onchip_memory_nios:readdata -> mm_interconnect_0:onchip_memory_nios_s1_readdata
	signal mm_interconnect_0_onchip_memory_nios_s1_address          : std_logic_vector(11 downto 0); -- mm_interconnect_0:onchip_memory_nios_s1_address -> onchip_memory_nios:address
	signal mm_interconnect_0_onchip_memory_nios_s1_byteenable       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory_nios_s1_byteenable -> onchip_memory_nios:byteenable
	signal mm_interconnect_0_onchip_memory_nios_s1_write            : std_logic;                     -- mm_interconnect_0:onchip_memory_nios_s1_write -> onchip_memory_nios:write
	signal mm_interconnect_0_onchip_memory_nios_s1_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory_nios_s1_writedata -> onchip_memory_nios:writedata
	signal mm_interconnect_0_onchip_memory_nios_s1_clken            : std_logic;                     -- mm_interconnect_0:onchip_memory_nios_s1_clken -> onchip_memory_nios:clken
	signal mm_interconnect_0_descriptor_memory_s1_chipselect        : std_logic;                     -- mm_interconnect_0:descriptor_memory_s1_chipselect -> descriptor_memory:chipselect
	signal mm_interconnect_0_descriptor_memory_s1_readdata          : std_logic_vector(31 downto 0); -- descriptor_memory:readdata -> mm_interconnect_0:descriptor_memory_s1_readdata
	signal mm_interconnect_0_descriptor_memory_s1_address           : std_logic_vector(9 downto 0);  -- mm_interconnect_0:descriptor_memory_s1_address -> descriptor_memory:address
	signal mm_interconnect_0_descriptor_memory_s1_byteenable        : std_logic_vector(3 downto 0);  -- mm_interconnect_0:descriptor_memory_s1_byteenable -> descriptor_memory:byteenable
	signal mm_interconnect_0_descriptor_memory_s1_write             : std_logic;                     -- mm_interconnect_0:descriptor_memory_s1_write -> descriptor_memory:write
	signal mm_interconnect_0_descriptor_memory_s1_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:descriptor_memory_s1_writedata -> descriptor_memory:writedata
	signal mm_interconnect_0_descriptor_memory_s1_clken             : std_logic;                     -- mm_interconnect_0:descriptor_memory_s1_clken -> descriptor_memory:clken
	signal irq_mapper_receiver0_irq                                 : std_logic;                     -- SGDMA_RX:csr_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                 : std_logic;                     -- SGDMA_TX:csr_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                 : std_logic;                     -- UART:av_irq -> irq_mapper:receiver2_irq
	signal nios2e_irq_irq                                           : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2e:irq
	signal demultiplexer_0_out0_valid                               : std_logic;                     -- demultiplexer_0:out0_valid -> avalon_st_adapter:in_0_valid
	signal demultiplexer_0_out0_data                                : std_logic_vector(31 downto 0); -- demultiplexer_0:out0_data -> avalon_st_adapter:in_0_data
	signal demultiplexer_0_out0_ready                               : std_logic;                     -- avalon_st_adapter:in_0_ready -> demultiplexer_0:out0_ready
	signal demultiplexer_0_out0_startofpacket                       : std_logic;                     -- demultiplexer_0:out0_startofpacket -> avalon_st_adapter:in_0_startofpacket
	signal demultiplexer_0_out0_endofpacket                         : std_logic;                     -- demultiplexer_0:out0_endofpacket -> avalon_st_adapter:in_0_endofpacket
	signal demultiplexer_0_out0_empty                               : std_logic_vector(1 downto 0);  -- demultiplexer_0:out0_empty -> avalon_st_adapter:in_0_empty
	signal avalon_st_adapter_out_0_valid                            : std_logic;                     -- avalon_st_adapter:out_0_valid -> SGDMA_RX:in_valid
	signal avalon_st_adapter_out_0_data                             : std_logic_vector(31 downto 0); -- avalon_st_adapter:out_0_data -> SGDMA_RX:in_data
	signal avalon_st_adapter_out_0_ready                            : std_logic;                     -- SGDMA_RX:in_ready -> avalon_st_adapter:out_0_ready
	signal avalon_st_adapter_out_0_startofpacket                    : std_logic;                     -- avalon_st_adapter:out_0_startofpacket -> SGDMA_RX:in_startofpacket
	signal avalon_st_adapter_out_0_endofpacket                      : std_logic;                     -- avalon_st_adapter:out_0_endofpacket -> SGDMA_RX:in_endofpacket
	signal avalon_st_adapter_out_0_error                            : std_logic_vector(5 downto 0);  -- avalon_st_adapter:out_0_error -> SGDMA_RX:in_error
	signal avalon_st_adapter_out_0_empty                            : std_logic_vector(1 downto 0);  -- avalon_st_adapter:out_0_empty -> SGDMA_RX:in_empty
	signal demultiplexer_0_out1_valid                               : std_logic;                     -- demultiplexer_0:out1_valid -> avalon_st_adapter_001:in_0_valid
	signal demultiplexer_0_out1_data                                : std_logic_vector(31 downto 0); -- demultiplexer_0:out1_data -> avalon_st_adapter_001:in_0_data
	signal demultiplexer_0_out1_ready                               : std_logic;                     -- avalon_st_adapter_001:in_0_ready -> demultiplexer_0:out1_ready
	signal demultiplexer_0_out1_startofpacket                       : std_logic;                     -- demultiplexer_0:out1_startofpacket -> avalon_st_adapter_001:in_0_startofpacket
	signal demultiplexer_0_out1_endofpacket                         : std_logic;                     -- demultiplexer_0:out1_endofpacket -> avalon_st_adapter_001:in_0_endofpacket
	signal demultiplexer_0_out1_empty                               : std_logic_vector(1 downto 0);  -- demultiplexer_0:out1_empty -> avalon_st_adapter_001:in_0_empty
	signal avalon_st_adapter_001_out_0_data                         : std_logic_vector(31 downto 0); -- avalon_st_adapter_001:out_0_data -> Filter_0:avsChannel
	signal avalon_st_adapter_001_out_0_startofpacket                : std_logic;                     -- avalon_st_adapter_001:out_0_startofpacket -> Filter_0:startofpacket
	signal avalon_st_adapter_001_out_0_endofpacket                  : std_logic;                     -- avalon_st_adapter_001:out_0_endofpacket -> Filter_0:endofpacket
	signal tse_mac_receive_valid                                    : std_logic;                     -- TSE_MAC:ff_rx_dval -> avalon_st_adapter_002:in_0_valid
	signal tse_mac_receive_data                                     : std_logic_vector(31 downto 0); -- TSE_MAC:ff_rx_data -> avalon_st_adapter_002:in_0_data
	signal tse_mac_receive_ready                                    : std_logic;                     -- avalon_st_adapter_002:in_0_ready -> TSE_MAC:ff_rx_rdy
	signal tse_mac_receive_startofpacket                            : std_logic;                     -- TSE_MAC:ff_rx_sop -> avalon_st_adapter_002:in_0_startofpacket
	signal tse_mac_receive_endofpacket                              : std_logic;                     -- TSE_MAC:ff_rx_eop -> avalon_st_adapter_002:in_0_endofpacket
	signal tse_mac_receive_error                                    : std_logic_vector(5 downto 0);  -- TSE_MAC:rx_err -> avalon_st_adapter_002:in_0_error
	signal tse_mac_receive_empty                                    : std_logic_vector(1 downto 0);  -- TSE_MAC:ff_rx_mod -> avalon_st_adapter_002:in_0_empty
	signal avalon_st_adapter_002_out_0_valid                        : std_logic;                     -- avalon_st_adapter_002:out_0_valid -> demultiplexer_0:in_valid
	signal avalon_st_adapter_002_out_0_data                         : std_logic_vector(31 downto 0); -- avalon_st_adapter_002:out_0_data -> demultiplexer_0:in_data
	signal avalon_st_adapter_002_out_0_ready                        : std_logic;                     -- demultiplexer_0:in_ready -> avalon_st_adapter_002:out_0_ready
	signal avalon_st_adapter_002_out_0_channel                      : std_logic;                     -- avalon_st_adapter_002:out_0_channel -> demultiplexer_0:in_channel
	signal avalon_st_adapter_002_out_0_startofpacket                : std_logic;                     -- avalon_st_adapter_002:out_0_startofpacket -> demultiplexer_0:in_startofpacket
	signal avalon_st_adapter_002_out_0_endofpacket                  : std_logic;                     -- avalon_st_adapter_002:out_0_endofpacket -> demultiplexer_0:in_endofpacket
	signal avalon_st_adapter_002_out_0_empty                        : std_logic_vector(1 downto 0);  -- avalon_st_adapter_002:out_0_empty -> demultiplexer_0:in_empty
	signal rst_controller_reset_out_reset                           : std_logic;                     -- rst_controller:reset_out -> [Filter_0:reset, TSE_MAC:reset, avalon_st_adapter_002:in_rst_0_reset, descriptor_memory:reset, irq_mapper:reset, mm_interconnect_0:nios2e_reset_reset_bridge_in_reset_reset, onchip_memory_nios:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                       : std_logic;                     -- rst_controller:reset_req -> [descriptor_memory:reset_req, nios2e:reset_req, onchip_memory_nios:reset_req, rst_translator:reset_req_in]
	signal rst_controller_001_reset_out_reset                       : std_logic;                     -- rst_controller_001:reset_out -> [avalon_st_adapter:in_rst_0_reset, avalon_st_adapter_001:in_rst_0_reset, rst_controller_001_reset_out_reset:in]
	signal mm_interconnect_0_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_uart_avalon_jtag_slave_read:inv -> UART:av_read_n
	signal mm_interconnect_0_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_uart_avalon_jtag_slave_write:inv -> UART:av_write_n
	signal rst_controller_reset_out_reset_ports_inv                 : std_logic;                     -- rst_controller_reset_out_reset:inv -> [SGDMA_RX:system_reset_n, SGDMA_TX:system_reset_n, UART:rst_n, nios2e:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv             : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> demultiplexer_0:reset_n

begin

	filter_0 : component PacketFilter
		port map (
			outData       => mm_interconnect_0_filter_0_avalon_slave_0_readdata,   --        avalon_slave_0.readdata
			inData        => mm_interconnect_0_filter_0_avalon_slave_0_writedata,  --                      .writedata
			address       => mm_interconnect_0_filter_0_avalon_slave_0_address,    --                      .address
			chipselect    => mm_interconnect_0_filter_0_avalon_slave_0_chipselect, --                      .chipselect
			readTo        => mm_interconnect_0_filter_0_avalon_slave_0_read,       --                      .read
			writeTo       => mm_interconnect_0_filter_0_avalon_slave_0_write,      --                      .write
			avsChannel    => avalon_st_adapter_001_out_0_data,                     -- avalon_streaming_sink.data
			startofpacket => avalon_st_adapter_001_out_0_startofpacket,            --                      .startofpacket
			endofpacket   => avalon_st_adapter_001_out_0_endofpacket,              --                      .endofpacket
			clock         => clk_clk,                                              --            clock_sink.clk
			reset         => rst_controller_reset_out_reset                        --            reset_sink.reset
		);

	sgdma_rx : component Wire_Shark_SGDMA_RX
		port map (
			clk                           => clk_clk,                                   --              clk.clk
			system_reset_n                => rst_controller_reset_out_reset_ports_inv,  --            reset.reset_n
			csr_chipselect                => mm_interconnect_0_sgdma_rx_csr_chipselect, --              csr.chipselect
			csr_address                   => mm_interconnect_0_sgdma_rx_csr_address,    --                 .address
			csr_read                      => mm_interconnect_0_sgdma_rx_csr_read,       --                 .read
			csr_write                     => mm_interconnect_0_sgdma_rx_csr_write,      --                 .write
			csr_writedata                 => mm_interconnect_0_sgdma_rx_csr_writedata,  --                 .writedata
			csr_readdata                  => mm_interconnect_0_sgdma_rx_csr_readdata,   --                 .readdata
			descriptor_read_readdata      => sgdma_rx_descriptor_read_readdata,         --  descriptor_read.readdata
			descriptor_read_readdatavalid => sgdma_rx_descriptor_read_readdatavalid,    --                 .readdatavalid
			descriptor_read_waitrequest   => sgdma_rx_descriptor_read_waitrequest,      --                 .waitrequest
			descriptor_read_address       => sgdma_rx_descriptor_read_address,          --                 .address
			descriptor_read_read          => sgdma_rx_descriptor_read_read,             --                 .read
			descriptor_write_waitrequest  => sgdma_rx_descriptor_write_waitrequest,     -- descriptor_write.waitrequest
			descriptor_write_address      => sgdma_rx_descriptor_write_address,         --                 .address
			descriptor_write_write        => sgdma_rx_descriptor_write_write,           --                 .write
			descriptor_write_writedata    => sgdma_rx_descriptor_write_writedata,       --                 .writedata
			csr_irq                       => irq_mapper_receiver0_irq,                  --          csr_irq.irq
			in_startofpacket              => avalon_st_adapter_out_0_startofpacket,     --               in.startofpacket
			in_endofpacket                => avalon_st_adapter_out_0_endofpacket,       --                 .endofpacket
			in_data                       => avalon_st_adapter_out_0_data,              --                 .data
			in_valid                      => avalon_st_adapter_out_0_valid,             --                 .valid
			in_ready                      => avalon_st_adapter_out_0_ready,             --                 .ready
			in_empty                      => avalon_st_adapter_out_0_empty,             --                 .empty
			in_error                      => avalon_st_adapter_out_0_error,             --                 .error
			m_write_waitrequest           => sgdma_rx_m_write_waitrequest,              --          m_write.waitrequest
			m_write_address               => sgdma_rx_m_write_address,                  --                 .address
			m_write_write                 => sgdma_rx_m_write_write,                    --                 .write
			m_write_writedata             => sgdma_rx_m_write_writedata,                --                 .writedata
			m_write_byteenable            => sgdma_rx_m_write_byteenable                --                 .byteenable
		);

	sgdma_tx : component Wire_Shark_SGDMA_TX
		port map (
			clk                           => clk_clk,                                   --              clk.clk
			system_reset_n                => rst_controller_reset_out_reset_ports_inv,  --            reset.reset_n
			csr_chipselect                => mm_interconnect_0_sgdma_tx_csr_chipselect, --              csr.chipselect
			csr_address                   => mm_interconnect_0_sgdma_tx_csr_address,    --                 .address
			csr_read                      => mm_interconnect_0_sgdma_tx_csr_read,       --                 .read
			csr_write                     => mm_interconnect_0_sgdma_tx_csr_write,      --                 .write
			csr_writedata                 => mm_interconnect_0_sgdma_tx_csr_writedata,  --                 .writedata
			csr_readdata                  => mm_interconnect_0_sgdma_tx_csr_readdata,   --                 .readdata
			descriptor_read_readdata      => sgdma_tx_descriptor_read_readdata,         --  descriptor_read.readdata
			descriptor_read_readdatavalid => sgdma_tx_descriptor_read_readdatavalid,    --                 .readdatavalid
			descriptor_read_waitrequest   => sgdma_tx_descriptor_read_waitrequest,      --                 .waitrequest
			descriptor_read_address       => sgdma_tx_descriptor_read_address,          --                 .address
			descriptor_read_read          => sgdma_tx_descriptor_read_read,             --                 .read
			descriptor_write_waitrequest  => sgdma_tx_descriptor_write_waitrequest,     -- descriptor_write.waitrequest
			descriptor_write_address      => sgdma_tx_descriptor_write_address,         --                 .address
			descriptor_write_write        => sgdma_tx_descriptor_write_write,           --                 .write
			descriptor_write_writedata    => sgdma_tx_descriptor_write_writedata,       --                 .writedata
			csr_irq                       => irq_mapper_receiver1_irq,                  --          csr_irq.irq
			m_read_readdata               => sgdma_tx_m_read_readdata,                  --           m_read.readdata
			m_read_readdatavalid          => sgdma_tx_m_read_readdatavalid,             --                 .readdatavalid
			m_read_waitrequest            => sgdma_tx_m_read_waitrequest,               --                 .waitrequest
			m_read_address                => sgdma_tx_m_read_address,                   --                 .address
			m_read_read                   => sgdma_tx_m_read_read,                      --                 .read
			out_data                      => sgdma_tx_out_data,                         --              out.data
			out_valid                     => sgdma_tx_out_valid,                        --                 .valid
			out_ready                     => sgdma_tx_out_ready,                        --                 .ready
			out_endofpacket               => sgdma_tx_out_endofpacket,                  --                 .endofpacket
			out_startofpacket             => sgdma_tx_out_startofpacket,                --                 .startofpacket
			out_empty                     => sgdma_tx_out_empty,                        --                 .empty
			out_error                     => sgdma_tx_out_error                         --                 .error
		);

	tse_mac : component Wire_Shark_TSE_MAC
		port map (
			clk           => clk_clk,                                            -- control_port_clock_connection.clk
			reset         => rst_controller_reset_out_reset,                     --              reset_connection.reset
			reg_addr      => mm_interconnect_0_tse_mac_control_port_address,     --                  control_port.address
			reg_data_out  => mm_interconnect_0_tse_mac_control_port_readdata,    --                              .readdata
			reg_rd        => mm_interconnect_0_tse_mac_control_port_read,        --                              .read
			reg_data_in   => mm_interconnect_0_tse_mac_control_port_writedata,   --                              .writedata
			reg_wr        => mm_interconnect_0_tse_mac_control_port_write,       --                              .write
			reg_busy      => mm_interconnect_0_tse_mac_control_port_waitrequest, --                              .waitrequest
			tx_clk        => pll_0_outclk0_clk,                                  --   pcs_mac_tx_clock_connection.clk
			rx_clk        => pll_0_outclk0_clk,                                  --   pcs_mac_rx_clock_connection.clk
			set_10        => eth_tse_0_mac_status_connection_set_10,             --         mac_status_connection.set_10
			set_1000      => eth_tse_0_mac_status_connection_set_1000,           --                              .set_1000
			eth_mode      => eth_tse_0_mac_status_connection_eth_mode,           --                              .eth_mode
			ena_10        => eth_tse_0_mac_status_connection_ena_10,             --                              .ena_10
			rgmii_in      => eth_tse_0_mac_rgmii_connection_rgmii_in,            --          mac_rgmii_connection.rgmii_in
			rgmii_out     => eth_tse_0_mac_rgmii_connection_rgmii_out,           --                              .rgmii_out
			rx_control    => eth_tse_0_mac_rgmii_connection_rx_control,          --                              .rx_control
			tx_control    => eth_tse_0_mac_rgmii_connection_tx_control,          --                              .tx_control
			ff_rx_clk     => clk_clk,                                            --      receive_clock_connection.clk
			ff_tx_clk     => clk_clk,                                            --     transmit_clock_connection.clk
			ff_rx_data    => tse_mac_receive_data,                               --                       receive.data
			ff_rx_eop     => tse_mac_receive_endofpacket,                        --                              .endofpacket
			rx_err        => tse_mac_receive_error,                              --                              .error
			ff_rx_mod     => tse_mac_receive_empty,                              --                              .empty
			ff_rx_rdy     => tse_mac_receive_ready,                              --                              .ready
			ff_rx_sop     => tse_mac_receive_startofpacket,                      --                              .startofpacket
			ff_rx_dval    => tse_mac_receive_valid,                              --                              .valid
			ff_tx_data    => sgdma_tx_out_data,                                  --                      transmit.data
			ff_tx_eop     => sgdma_tx_out_endofpacket,                           --                              .endofpacket
			ff_tx_err     => sgdma_tx_out_error,                                 --                              .error
			ff_tx_mod     => sgdma_tx_out_empty,                                 --                              .empty
			ff_tx_rdy     => sgdma_tx_out_ready,                                 --                              .ready
			ff_tx_sop     => sgdma_tx_out_startofpacket,                         --                              .startofpacket
			ff_tx_wren    => sgdma_tx_out_valid,                                 --                              .valid
			mdc           => eth_tse_0_mac_mdio_connection_mdc,                  --           mac_mdio_connection.mdc
			mdio_in       => eth_tse_0_mac_mdio_connection_mdio_in,              --                              .mdio_in
			mdio_out      => eth_tse_0_mac_mdio_connection_mdio_out,             --                              .mdio_out
			mdio_oen      => eth_tse_0_mac_mdio_connection_mdio_oen,             --                              .mdio_oen
			magic_wakeup  => open,                                               --           mac_misc_connection.magic_wakeup
			magic_sleep_n => open,                                               --                              .magic_sleep_n
			ff_tx_crc_fwd => open,                                               --                              .ff_tx_crc_fwd
			ff_tx_septy   => open,                                               --                              .ff_tx_septy
			tx_ff_uflow   => open,                                               --                              .tx_ff_uflow
			ff_tx_a_full  => open,                                               --                              .ff_tx_a_full
			ff_tx_a_empty => open,                                               --                              .ff_tx_a_empty
			rx_err_stat   => open,                                               --                              .rx_err_stat
			rx_frm_type   => open,                                               --                              .rx_frm_type
			ff_rx_dsav    => open,                                               --                              .ff_rx_dsav
			ff_rx_a_full  => open,                                               --                              .ff_rx_a_full
			ff_rx_a_empty => open                                                --                              .ff_rx_a_empty
		);

	uart : component Wire_Shark_UART
		port map (
			clk            => clk_clk,                                                  --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                 --             reset.reset_n
			av_chipselect  => mm_interconnect_0_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver2_irq                                  --               irq.irq
		);

	demultiplexer_0 : component Wire_Shark_demultiplexer_0
		port map (
			clk                => clk_clk,                                      --   clk.clk
			reset_n            => rst_controller_001_reset_out_reset_ports_inv, -- reset.reset_n
			in_data            => avalon_st_adapter_002_out_0_data,             --    in.data
			in_valid           => avalon_st_adapter_002_out_0_valid,            --      .valid
			in_ready           => avalon_st_adapter_002_out_0_ready,            --      .ready
			in_startofpacket   => avalon_st_adapter_002_out_0_startofpacket,    --      .startofpacket
			in_endofpacket     => avalon_st_adapter_002_out_0_endofpacket,      --      .endofpacket
			in_empty           => avalon_st_adapter_002_out_0_empty,            --      .empty
			in_channel         => avalon_st_adapter_002_out_0_channel,          --      .channel
			out0_data          => demultiplexer_0_out0_data,                    --  out0.data
			out0_valid         => demultiplexer_0_out0_valid,                   --      .valid
			out0_ready         => demultiplexer_0_out0_ready,                   --      .ready
			out0_startofpacket => demultiplexer_0_out0_startofpacket,           --      .startofpacket
			out0_endofpacket   => demultiplexer_0_out0_endofpacket,             --      .endofpacket
			out0_empty         => demultiplexer_0_out0_empty,                   --      .empty
			out1_data          => demultiplexer_0_out1_data,                    --  out1.data
			out1_valid         => demultiplexer_0_out1_valid,                   --      .valid
			out1_ready         => demultiplexer_0_out1_ready,                   --      .ready
			out1_startofpacket => demultiplexer_0_out1_startofpacket,           --      .startofpacket
			out1_endofpacket   => demultiplexer_0_out1_endofpacket,             --      .endofpacket
			out1_empty         => demultiplexer_0_out1_empty                    --      .empty
		);

	descriptor_memory : component Wire_Shark_descriptor_memory
		port map (
			clk        => clk_clk,                                           --   clk1.clk
			address    => mm_interconnect_0_descriptor_memory_s1_address,    --     s1.address
			clken      => mm_interconnect_0_descriptor_memory_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_descriptor_memory_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_descriptor_memory_s1_write,      --       .write
			readdata   => mm_interconnect_0_descriptor_memory_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_descriptor_memory_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_descriptor_memory_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                    -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,                --       .reset_req
			freeze     => '0'                                                -- (terminated)
		);

	nios2e : component Wire_Shark_nios2e
		port map (
			clk                                 => clk_clk,                                              --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,             --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                   --                          .reset_req
			d_address                           => nios2e_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2e_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2e_data_master_read,                              --                          .read
			d_readdata                          => nios2e_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2e_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2e_data_master_write,                             --                          .write
			d_writedata                         => nios2e_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2e_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2e_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2e_instruction_master_read,                       --                          .read
			i_readdata                          => nios2e_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2e_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios2e_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2e_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2e_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2e_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2e_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2e_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2e_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2e_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2e_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2e_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                  -- custom_instruction_master.readra
		);

	onchip_memory_nios : component Wire_Shark_onchip_memory_nios
		port map (
			clk        => clk_clk,                                            --   clk1.clk
			address    => mm_interconnect_0_onchip_memory_nios_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory_nios_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory_nios_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory_nios_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory_nios_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory_nios_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory_nios_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                     -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,                 --       .reset_req
			freeze     => '0'                                                 -- (terminated)
		);

	pll_0 : component Wire_Shark_pll_0
		port map (
			refclk   => clk_clk,                          --  refclk.clk
			rst      => nios2e_debug_reset_request_reset, --   reset.reset
			outclk_0 => pll_0_outclk0_clk,                -- outclk0.clk
			locked   => open                              --  locked.export
		);

	mm_interconnect_0 : component Wire_Shark_mm_interconnect_0
		port map (
			clk_0_clk_clk                            => clk_clk,                                              --                          clk_0_clk.clk
			nios2e_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                       -- nios2e_reset_reset_bridge_in_reset.reset
			nios2e_data_master_address               => nios2e_data_master_address,                           --                 nios2e_data_master.address
			nios2e_data_master_waitrequest           => nios2e_data_master_waitrequest,                       --                                   .waitrequest
			nios2e_data_master_byteenable            => nios2e_data_master_byteenable,                        --                                   .byteenable
			nios2e_data_master_read                  => nios2e_data_master_read,                              --                                   .read
			nios2e_data_master_readdata              => nios2e_data_master_readdata,                          --                                   .readdata
			nios2e_data_master_write                 => nios2e_data_master_write,                             --                                   .write
			nios2e_data_master_writedata             => nios2e_data_master_writedata,                         --                                   .writedata
			nios2e_data_master_debugaccess           => nios2e_data_master_debugaccess,                       --                                   .debugaccess
			nios2e_instruction_master_address        => nios2e_instruction_master_address,                    --          nios2e_instruction_master.address
			nios2e_instruction_master_waitrequest    => nios2e_instruction_master_waitrequest,                --                                   .waitrequest
			nios2e_instruction_master_read           => nios2e_instruction_master_read,                       --                                   .read
			nios2e_instruction_master_readdata       => nios2e_instruction_master_readdata,                   --                                   .readdata
			SGDMA_RX_descriptor_read_address         => sgdma_rx_descriptor_read_address,                     --           SGDMA_RX_descriptor_read.address
			SGDMA_RX_descriptor_read_waitrequest     => sgdma_rx_descriptor_read_waitrequest,                 --                                   .waitrequest
			SGDMA_RX_descriptor_read_read            => sgdma_rx_descriptor_read_read,                        --                                   .read
			SGDMA_RX_descriptor_read_readdata        => sgdma_rx_descriptor_read_readdata,                    --                                   .readdata
			SGDMA_RX_descriptor_read_readdatavalid   => sgdma_rx_descriptor_read_readdatavalid,               --                                   .readdatavalid
			SGDMA_RX_descriptor_write_address        => sgdma_rx_descriptor_write_address,                    --          SGDMA_RX_descriptor_write.address
			SGDMA_RX_descriptor_write_waitrequest    => sgdma_rx_descriptor_write_waitrequest,                --                                   .waitrequest
			SGDMA_RX_descriptor_write_write          => sgdma_rx_descriptor_write_write,                      --                                   .write
			SGDMA_RX_descriptor_write_writedata      => sgdma_rx_descriptor_write_writedata,                  --                                   .writedata
			SGDMA_RX_m_write_address                 => sgdma_rx_m_write_address,                             --                   SGDMA_RX_m_write.address
			SGDMA_RX_m_write_waitrequest             => sgdma_rx_m_write_waitrequest,                         --                                   .waitrequest
			SGDMA_RX_m_write_byteenable              => sgdma_rx_m_write_byteenable,                          --                                   .byteenable
			SGDMA_RX_m_write_write                   => sgdma_rx_m_write_write,                               --                                   .write
			SGDMA_RX_m_write_writedata               => sgdma_rx_m_write_writedata,                           --                                   .writedata
			SGDMA_TX_descriptor_read_address         => sgdma_tx_descriptor_read_address,                     --           SGDMA_TX_descriptor_read.address
			SGDMA_TX_descriptor_read_waitrequest     => sgdma_tx_descriptor_read_waitrequest,                 --                                   .waitrequest
			SGDMA_TX_descriptor_read_read            => sgdma_tx_descriptor_read_read,                        --                                   .read
			SGDMA_TX_descriptor_read_readdata        => sgdma_tx_descriptor_read_readdata,                    --                                   .readdata
			SGDMA_TX_descriptor_read_readdatavalid   => sgdma_tx_descriptor_read_readdatavalid,               --                                   .readdatavalid
			SGDMA_TX_descriptor_write_address        => sgdma_tx_descriptor_write_address,                    --          SGDMA_TX_descriptor_write.address
			SGDMA_TX_descriptor_write_waitrequest    => sgdma_tx_descriptor_write_waitrequest,                --                                   .waitrequest
			SGDMA_TX_descriptor_write_write          => sgdma_tx_descriptor_write_write,                      --                                   .write
			SGDMA_TX_descriptor_write_writedata      => sgdma_tx_descriptor_write_writedata,                  --                                   .writedata
			SGDMA_TX_m_read_address                  => sgdma_tx_m_read_address,                              --                    SGDMA_TX_m_read.address
			SGDMA_TX_m_read_waitrequest              => sgdma_tx_m_read_waitrequest,                          --                                   .waitrequest
			SGDMA_TX_m_read_read                     => sgdma_tx_m_read_read,                                 --                                   .read
			SGDMA_TX_m_read_readdata                 => sgdma_tx_m_read_readdata,                             --                                   .readdata
			SGDMA_TX_m_read_readdatavalid            => sgdma_tx_m_read_readdatavalid,                        --                                   .readdatavalid
			descriptor_memory_s1_address             => mm_interconnect_0_descriptor_memory_s1_address,       --               descriptor_memory_s1.address
			descriptor_memory_s1_write               => mm_interconnect_0_descriptor_memory_s1_write,         --                                   .write
			descriptor_memory_s1_readdata            => mm_interconnect_0_descriptor_memory_s1_readdata,      --                                   .readdata
			descriptor_memory_s1_writedata           => mm_interconnect_0_descriptor_memory_s1_writedata,     --                                   .writedata
			descriptor_memory_s1_byteenable          => mm_interconnect_0_descriptor_memory_s1_byteenable,    --                                   .byteenable
			descriptor_memory_s1_chipselect          => mm_interconnect_0_descriptor_memory_s1_chipselect,    --                                   .chipselect
			descriptor_memory_s1_clken               => mm_interconnect_0_descriptor_memory_s1_clken,         --                                   .clken
			Filter_0_avalon_slave_0_address          => mm_interconnect_0_filter_0_avalon_slave_0_address,    --            Filter_0_avalon_slave_0.address
			Filter_0_avalon_slave_0_write            => mm_interconnect_0_filter_0_avalon_slave_0_write,      --                                   .write
			Filter_0_avalon_slave_0_read             => mm_interconnect_0_filter_0_avalon_slave_0_read,       --                                   .read
			Filter_0_avalon_slave_0_readdata         => mm_interconnect_0_filter_0_avalon_slave_0_readdata,   --                                   .readdata
			Filter_0_avalon_slave_0_writedata        => mm_interconnect_0_filter_0_avalon_slave_0_writedata,  --                                   .writedata
			Filter_0_avalon_slave_0_chipselect       => mm_interconnect_0_filter_0_avalon_slave_0_chipselect, --                                   .chipselect
			nios2e_debug_mem_slave_address           => mm_interconnect_0_nios2e_debug_mem_slave_address,     --             nios2e_debug_mem_slave.address
			nios2e_debug_mem_slave_write             => mm_interconnect_0_nios2e_debug_mem_slave_write,       --                                   .write
			nios2e_debug_mem_slave_read              => mm_interconnect_0_nios2e_debug_mem_slave_read,        --                                   .read
			nios2e_debug_mem_slave_readdata          => mm_interconnect_0_nios2e_debug_mem_slave_readdata,    --                                   .readdata
			nios2e_debug_mem_slave_writedata         => mm_interconnect_0_nios2e_debug_mem_slave_writedata,   --                                   .writedata
			nios2e_debug_mem_slave_byteenable        => mm_interconnect_0_nios2e_debug_mem_slave_byteenable,  --                                   .byteenable
			nios2e_debug_mem_slave_waitrequest       => mm_interconnect_0_nios2e_debug_mem_slave_waitrequest, --                                   .waitrequest
			nios2e_debug_mem_slave_debugaccess       => mm_interconnect_0_nios2e_debug_mem_slave_debugaccess, --                                   .debugaccess
			onchip_memory_nios_s1_address            => mm_interconnect_0_onchip_memory_nios_s1_address,      --              onchip_memory_nios_s1.address
			onchip_memory_nios_s1_write              => mm_interconnect_0_onchip_memory_nios_s1_write,        --                                   .write
			onchip_memory_nios_s1_readdata           => mm_interconnect_0_onchip_memory_nios_s1_readdata,     --                                   .readdata
			onchip_memory_nios_s1_writedata          => mm_interconnect_0_onchip_memory_nios_s1_writedata,    --                                   .writedata
			onchip_memory_nios_s1_byteenable         => mm_interconnect_0_onchip_memory_nios_s1_byteenable,   --                                   .byteenable
			onchip_memory_nios_s1_chipselect         => mm_interconnect_0_onchip_memory_nios_s1_chipselect,   --                                   .chipselect
			onchip_memory_nios_s1_clken              => mm_interconnect_0_onchip_memory_nios_s1_clken,        --                                   .clken
			SGDMA_RX_csr_address                     => mm_interconnect_0_sgdma_rx_csr_address,               --                       SGDMA_RX_csr.address
			SGDMA_RX_csr_write                       => mm_interconnect_0_sgdma_rx_csr_write,                 --                                   .write
			SGDMA_RX_csr_read                        => mm_interconnect_0_sgdma_rx_csr_read,                  --                                   .read
			SGDMA_RX_csr_readdata                    => mm_interconnect_0_sgdma_rx_csr_readdata,              --                                   .readdata
			SGDMA_RX_csr_writedata                   => mm_interconnect_0_sgdma_rx_csr_writedata,             --                                   .writedata
			SGDMA_RX_csr_chipselect                  => mm_interconnect_0_sgdma_rx_csr_chipselect,            --                                   .chipselect
			SGDMA_TX_csr_address                     => mm_interconnect_0_sgdma_tx_csr_address,               --                       SGDMA_TX_csr.address
			SGDMA_TX_csr_write                       => mm_interconnect_0_sgdma_tx_csr_write,                 --                                   .write
			SGDMA_TX_csr_read                        => mm_interconnect_0_sgdma_tx_csr_read,                  --                                   .read
			SGDMA_TX_csr_readdata                    => mm_interconnect_0_sgdma_tx_csr_readdata,              --                                   .readdata
			SGDMA_TX_csr_writedata                   => mm_interconnect_0_sgdma_tx_csr_writedata,             --                                   .writedata
			SGDMA_TX_csr_chipselect                  => mm_interconnect_0_sgdma_tx_csr_chipselect,            --                                   .chipselect
			TSE_MAC_control_port_address             => mm_interconnect_0_tse_mac_control_port_address,       --               TSE_MAC_control_port.address
			TSE_MAC_control_port_write               => mm_interconnect_0_tse_mac_control_port_write,         --                                   .write
			TSE_MAC_control_port_read                => mm_interconnect_0_tse_mac_control_port_read,          --                                   .read
			TSE_MAC_control_port_readdata            => mm_interconnect_0_tse_mac_control_port_readdata,      --                                   .readdata
			TSE_MAC_control_port_writedata           => mm_interconnect_0_tse_mac_control_port_writedata,     --                                   .writedata
			TSE_MAC_control_port_waitrequest         => mm_interconnect_0_tse_mac_control_port_waitrequest,   --                                   .waitrequest
			UART_avalon_jtag_slave_address           => mm_interconnect_0_uart_avalon_jtag_slave_address,     --             UART_avalon_jtag_slave.address
			UART_avalon_jtag_slave_write             => mm_interconnect_0_uart_avalon_jtag_slave_write,       --                                   .write
			UART_avalon_jtag_slave_read              => mm_interconnect_0_uart_avalon_jtag_slave_read,        --                                   .read
			UART_avalon_jtag_slave_readdata          => mm_interconnect_0_uart_avalon_jtag_slave_readdata,    --                                   .readdata
			UART_avalon_jtag_slave_writedata         => mm_interconnect_0_uart_avalon_jtag_slave_writedata,   --                                   .writedata
			UART_avalon_jtag_slave_waitrequest       => mm_interconnect_0_uart_avalon_jtag_slave_waitrequest, --                                   .waitrequest
			UART_avalon_jtag_slave_chipselect        => mm_interconnect_0_uart_avalon_jtag_slave_chipselect   --                                   .chipselect
		);

	irq_mapper : component Wire_Shark_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			sender_irq    => nios2e_irq_irq                  --    sender.irq
		);

	avalon_st_adapter : component Wire_Shark_avalon_st_adapter
		generic map (
			inBitsPerSymbol => 8,
			inUsePackets    => 1,
			inDataWidth     => 32,
			inChannelWidth  => 0,
			inErrorWidth    => 0,
			inUseEmptyPort  => 1,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 0,
			outDataWidth    => 32,
			outChannelWidth => 0,
			outErrorWidth   => 6,
			outUseEmptyPort => 1,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk        => clk_clk,                               -- in_clk_0.clk
			in_rst_0_reset      => rst_controller_001_reset_out_reset,    -- in_rst_0.reset
			in_0_data           => demultiplexer_0_out0_data,             --     in_0.data
			in_0_valid          => demultiplexer_0_out0_valid,            --         .valid
			in_0_ready          => demultiplexer_0_out0_ready,            --         .ready
			in_0_startofpacket  => demultiplexer_0_out0_startofpacket,    --         .startofpacket
			in_0_endofpacket    => demultiplexer_0_out0_endofpacket,      --         .endofpacket
			in_0_empty          => demultiplexer_0_out0_empty,            --         .empty
			out_0_data          => avalon_st_adapter_out_0_data,          --    out_0.data
			out_0_valid         => avalon_st_adapter_out_0_valid,         --         .valid
			out_0_ready         => avalon_st_adapter_out_0_ready,         --         .ready
			out_0_startofpacket => avalon_st_adapter_out_0_startofpacket, --         .startofpacket
			out_0_endofpacket   => avalon_st_adapter_out_0_endofpacket,   --         .endofpacket
			out_0_empty         => avalon_st_adapter_out_0_empty,         --         .empty
			out_0_error         => avalon_st_adapter_out_0_error          --         .error
		);

	avalon_st_adapter_001 : component Wire_Shark_avalon_st_adapter_001
		generic map (
			inBitsPerSymbol => 8,
			inUsePackets    => 1,
			inDataWidth     => 32,
			inChannelWidth  => 0,
			inErrorWidth    => 0,
			inUseEmptyPort  => 1,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 0,
			outDataWidth    => 32,
			outChannelWidth => 0,
			outErrorWidth   => 0,
			outUseEmptyPort => 0,
			outUseValid     => 0,
			outUseReady     => 0,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk        => clk_clk,                                   -- in_clk_0.clk
			in_rst_0_reset      => rst_controller_001_reset_out_reset,        -- in_rst_0.reset
			in_0_data           => demultiplexer_0_out1_data,                 --     in_0.data
			in_0_valid          => demultiplexer_0_out1_valid,                --         .valid
			in_0_ready          => demultiplexer_0_out1_ready,                --         .ready
			in_0_startofpacket  => demultiplexer_0_out1_startofpacket,        --         .startofpacket
			in_0_endofpacket    => demultiplexer_0_out1_endofpacket,          --         .endofpacket
			in_0_empty          => demultiplexer_0_out1_empty,                --         .empty
			out_0_data          => avalon_st_adapter_001_out_0_data,          --    out_0.data
			out_0_startofpacket => avalon_st_adapter_001_out_0_startofpacket, --         .startofpacket
			out_0_endofpacket   => avalon_st_adapter_001_out_0_endofpacket    --         .endofpacket
		);

	avalon_st_adapter_002 : component Wire_Shark_avalon_st_adapter_002
		generic map (
			inBitsPerSymbol => 8,
			inUsePackets    => 1,
			inDataWidth     => 32,
			inChannelWidth  => 0,
			inErrorWidth    => 6,
			inUseEmptyPort  => 1,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 2,
			outDataWidth    => 32,
			outChannelWidth => 1,
			outErrorWidth   => 0,
			outUseEmptyPort => 1,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk        => clk_clk,                                   -- in_clk_0.clk
			in_rst_0_reset      => rst_controller_reset_out_reset,            -- in_rst_0.reset
			in_0_data           => tse_mac_receive_data,                      --     in_0.data
			in_0_valid          => tse_mac_receive_valid,                     --         .valid
			in_0_ready          => tse_mac_receive_ready,                     --         .ready
			in_0_startofpacket  => tse_mac_receive_startofpacket,             --         .startofpacket
			in_0_endofpacket    => tse_mac_receive_endofpacket,               --         .endofpacket
			in_0_empty          => tse_mac_receive_empty,                     --         .empty
			in_0_error          => tse_mac_receive_error,                     --         .error
			out_0_data          => avalon_st_adapter_002_out_0_data,          --    out_0.data
			out_0_valid         => avalon_st_adapter_002_out_0_valid,         --         .valid
			out_0_ready         => avalon_st_adapter_002_out_0_ready,         --         .ready
			out_0_startofpacket => avalon_st_adapter_002_out_0_startofpacket, --         .startofpacket
			out_0_endofpacket   => avalon_st_adapter_002_out_0_endofpacket,   --         .endofpacket
			out_0_empty         => avalon_st_adapter_002_out_0_empty,         --         .empty
			out_0_channel       => avalon_st_adapter_002_out_0_channel        --         .channel
		);

	rst_controller : component wire_shark_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2e_debug_reset_request_reset,   -- reset_in0.reset
			reset_in1      => nios2e_debug_reset_request_reset,   -- reset_in1.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component wire_shark_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2e_debug_reset_request_reset,   -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	mm_interconnect_0_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_uart_avalon_jtag_slave_read;

	mm_interconnect_0_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_uart_avalon_jtag_slave_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of Wire_Shark
